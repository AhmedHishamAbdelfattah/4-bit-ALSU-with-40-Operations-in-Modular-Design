module ALSU_Top_Module_TB ;

  parameter Width = 4; 
  parameter Width_Sel = 6;          
  parameter Output_Width = 4;    
  parameter Delay = 10;    

  reg [Width-1:0] A , B ; 
  reg [Width_Sel-1:0] Sel ;
  wire [Output_Width-1:0] Out ;
  wire carry_out ;
  wire Negative_Sign_Flag ;
  integer error_count = 0;

ALSU_Top_Module DUT ( .A ( A ) ,
                      .B ( B ) , 
                      .Sel ( Sel ) ,
                      .Out ( Out ) ,
                      .Carry_Out ( carry_out ) ,
                      .Negative_Sign_Flag( Negative_Sign_Flag )
                    );

  initial begin
  $monitor("A = %b , B = %b , Sel = %b , Out = %b , Carry_Out = %b , Negative_Sign_Flag = %b" ,
            A , B , Sel , Out , Out , carry_out , Negative_Sign_Flag);
  end
  
  initial begin 
// -------------------------------------------------------------------------------------------------------------------------------

// Arithmetic & Arithmetical Shift Operations

  // when Sel is 6'b000000 which indicates A + B 
  run_test(4'b0101, 4'b0100, 6'b000000, 4'b1001, 1'b0, 1'b0); // 5 + 4 = 9
  run_test(4'b0101, 4'b0011, 6'b000000, 4'b1000, 1'b0, 1'b0); // 5 + 3 = 8
  run_test(4'b0000, 4'b0000, 6'b000000, 4'b0000, 1'b0, 1'b0); // 0 + 0 = 0
  run_test(4'b1111, 4'b0011, 6'b000000, 4'b0010, 1'b1, 1'b0); // 15 + 3 = 18 → 0010 + carry
  run_test(4'b0011, 4'b0101, 6'b000000, 4'b1000, 1'b0, 1'b0); // 3 + 5 = 8
  run_test(4'b1010, 4'b0001, 6'b000000, 4'b1011, 1'b0, 1'b0); // 10 + 1 = 11
  run_test(4'b1100, 4'b1101, 6'b000000, 4'b1001, 1'b1, 1'b0); // 12 + 13 = 25 → 1001 + carry

  // when Sel is 6'b000001 which indicates A - B 
  run_test(4'b0101, 4'b0100, 6'b000001, 4'b0001, 1'b0, 1'b0); // 5 - 4 = 1
  run_test(4'b0101, 4'b0011, 6'b000001, 4'b0010, 1'b0, 1'b0); // 5 - 3 = 2
  run_test(4'b0000, 4'b0000, 6'b000001, 4'b0000, 1'b0, 1'b0); // 0 - 0 = 0
  run_test(4'b1111, 4'b0011, 6'b000001, 4'b1100, 1'b0, 1'b0); // 15 - 3 = 12 → 1100
  run_test(4'b0011, 4'b0101, 6'b000001, 4'b1110, 1'b0, 1'b1); // 3 - 5 = -2 → 0010 (negative)
  run_test(4'b1010, 4'b0001, 6'b000001, 4'b1001, 1'b0, 1'b0); // 10 - 1 = 9
  run_test(4'b1100, 4'b1101, 6'b000001, 4'b1111, 1'b0, 1'b1); // 12 - 13 = -1 → 0001 (negative)

  // when Sel is 6'b000010 which indicates 2's Comp.(B)
  run_test(4'b0101, 4'b1100, 6'b000010, 4'b0100, 1'b0, 1'b0); // ~1100+1 = 0011+1 = 0100
  run_test(4'b0101, 4'b0101, 6'b000010, 4'b1011, 1'b0, 1'b0); // ~0101+1 = 1010+1 = 1011
  run_test(4'b0101, 4'b1111, 6'b000010, 4'b0001, 1'b0, 1'b0); // ~1111+1 = 0000+1 = 0001
  run_test(4'b0101, 4'b0011, 6'b000010, 4'b1101, 1'b0, 1'b0); // ~0011+1 = 1100+1 = 1101
  run_test(4'b0101, 4'b1010, 6'b000010, 4'b0110, 1'b0, 1'b0); // ~1010+1 = 0101+1 = 0110
  run_test(4'b0101, 4'b1101, 6'b000010, 4'b0011, 1'b0, 1'b0); // ~1101+1 = 0010+1 = 0011
  run_test(4'b0101, 4'b0001, 6'b000010, 4'b1111, 1'b0, 1'b0); // ~0001+1 = 1110+1 = 1111
  run_test(4'b0101, 4'b0010, 6'b000010, 4'b1110, 1'b0, 1'b0); // ~0010+1 = 1101+1 = 1110
  run_test(4'b0101, 4'b1000, 6'b000010, 4'b1000, 1'b0, 1'b0); // ~1000+1 = 0111+1 = 1000 

  // when Sel is 6'b000011 which indicates 2's Comp.(A)
  run_test(4'b0101, 4'b1000, 6'b000011, 4'b1011, 1'b0, 1'b0); // ~0101+1 = 1010+1 = 1011
  run_test(4'b1100, 4'b1000, 6'b000011, 4'b0100, 1'b0, 1'b0); // ~1100+1 = 0011+1 = 0100
  run_test(4'b0001, 4'b1000, 6'b000011, 4'b1111, 1'b0, 1'b0); // ~0001+1 = 1110+1 = 1111
  run_test(4'b0011, 4'b1000, 6'b000011, 4'b1101, 1'b0, 1'b0); // ~0011+1 = 1100+1 = 1101
  run_test(4'b1010, 4'b1000, 6'b000011, 4'b0110, 1'b0, 1'b0); // ~1010+1 = 0101+1 = 0110
  run_test(4'b1101, 4'b1000, 6'b000011, 4'b0011, 1'b0, 1'b0); // ~1101+1 = 0010+1 = 0011
  run_test(4'b0010, 4'b1000, 6'b000011, 4'b1110, 1'b0, 1'b0); // ~0010+1 = 1101+1 = 1110
  run_test(4'b1000, 4'b1000, 6'b000011, 4'b1000, 1'b0, 1'b0); // ~1000+1 = 0111+1 = 1000


  // when Sel is 6'b000100 which indicates A * B ( Least Significant 4-bits )
  run_test(4'b0101, 4'b1000, 6'b000100, 4'b1000, 1'b0, 1'b0); // 5*8 = 40 → 00101000 → LSB = 1000
  run_test(4'b1100, 4'b1000, 6'b000100, 4'b0000, 1'b0, 1'b0); // 12*8 = 96 → 01100000 → LSB = 0000
  run_test(4'b0001, 4'b1000, 6'b000100, 4'b1000, 1'b0, 1'b0); // 1*8 = 8 → 00001000 → LSB = 1000 
  run_test(4'b0011, 4'b1000, 6'b000100, 4'b1000, 1'b0, 1'b0); // 3*8 = 24 → 00011000 → LSB = 1000 
  run_test(4'b1010, 4'b1000, 6'b000100, 4'b0000, 1'b0, 1'b0); // 10*8 = 80 → 01010000 → LSB = 0000
  run_test(4'b1101, 4'b1000, 6'b000100, 4'b1000, 1'b0, 1'b0); // 13*8 = 104 → 01101000 → LSB = 1000
  run_test(4'b0001, 4'b0011, 6'b000100, 4'b0011, 1'b0, 1'b0); // 1*3 = 3 → 00000011 → LSB = 0011
  run_test(4'b0010, 4'b0101, 6'b000100, 4'b1010, 1'b0, 1'b0); // 2*5 = 10 → 00001010 → LSB = 1010
  run_test(4'b1111, 4'b1111, 6'b000100, 4'b0001, 1'b0, 1'b0); // 15*15 = 11100001 →  → LSB = 0001

  // when Sel is 6'b000101 which indicates A * B ( Most Significant 4-bits ) 
  run_test(4'b0101, 4'b1000, 6'b000101, 4'b0010, 1'b0, 1'b0); // 5*8 = 40 → 00101000 → MSB = 0010
  run_test(4'b1100, 4'b1000, 6'b000101, 4'b0110, 1'b0, 1'b0); // 12*8 = 96 → 01100000 → MSB = 0110
  run_test(4'b0001, 4'b1000, 6'b000101, 4'b0000, 1'b0, 1'b0); // 1*8 = 8 → 00001000 → MSB = 0000  
  run_test(4'b0011, 4'b1000, 6'b000101, 4'b0001, 1'b0, 1'b0); // 3*8 = 24 → 00011000 → MSB = 0001 
  run_test(4'b1010, 4'b1000, 6'b000101, 4'b0101, 1'b0, 1'b0); // 10*8 = 80 → 01010000 → MSB = 0101
  run_test(4'b1101, 4'b1000, 6'b000101, 4'b0110, 1'b0, 1'b0); // 13*8 = 104 → 01101000 → MSB = 0110
  run_test(4'b0001, 4'b0011, 6'b000101, 4'b0000, 1'b0, 1'b0); // 1*3 = 3 → 00000011 → MSB = 0000
  run_test(4'b0010, 4'b0101, 6'b000101, 4'b0000, 1'b0, 1'b0); // 2*5 = 10 → 00001010 → MSB = 0000
  run_test(4'b1111, 4'b1111, 6'b000101, 4'b1110, 1'b0, 1'b0); // 15*15 = 11100001 →  → MSB = 1110

  // when Sel is 6'b001100 which indicates A / B ( Quotient ) 
  run_test(4'b0101, 4'b0010, 6'b001100, 4'b0010, 1'b0, 1'b0); // 5 / 2 = 2
  run_test(4'b1100, 4'b0011, 6'b001100, 4'b0100, 1'b0, 1'b0); // 12 / 3 = 4
  run_test(4'b0110, 4'b0011, 6'b001100, 4'b0010, 1'b0, 1'b0); // 6 / 3 = 2
  run_test(4'b1010, 4'b0100, 6'b001100, 4'b0010, 1'b0, 1'b0); // 10 / 4 = 2
  run_test(4'b1110, 4'b0101, 6'b001100, 4'b0010, 1'b0, 1'b0); // 14 / 5 = 2
  run_test(4'b0111, 4'b0010, 6'b001100, 4'b0011, 1'b0, 1'b0); // 7 / 2 = 3
  run_test(4'b1000, 4'b0100, 6'b001100, 4'b0010, 1'b0, 1'b0); // 8 / 4 = 2
  run_test(4'b0010, 4'b0101, 6'b001100, 4'b0000, 1'b0, 1'b0); // 2 / 5 = 0
  run_test(4'b1000, 4'b0011, 6'b001100, 4'b0010, 1'b0, 1'b0); // 8 / 3 = 2

  // when Sel is 6'b001101 which indicates A / B ( Remainder ) 
  run_test(4'b0101, 4'b0010, 6'b001101, 4'b0001, 1'b0, 1'b0); // 5 % 2 = 1
  run_test(4'b1100, 4'b0011, 6'b001101, 4'b0000, 1'b0, 1'b0); // 12 % 3 = 0
  run_test(4'b0110, 4'b0011, 6'b001101, 4'b0000, 1'b0, 1'b0); // 6 % 3 = 0
  run_test(4'b1010, 4'b0100, 6'b001101, 4'b0010, 1'b0, 1'b0); // 10 % 4 = 2
  run_test(4'b1110, 4'b0101, 6'b001101, 4'b0000, 1'b0, 1'b0); // 14 % 5 = 4
  run_test(4'b0111, 4'b0010, 6'b001101, 4'b0001, 1'b0, 1'b0); // 7 % 2 = 1
  run_test(4'b1000, 4'b0100, 6'b001101, 4'b0000, 1'b0, 1'b0); // 8 % 4 = 0
  run_test(4'b0010, 4'b0101, 6'b001101, 4'b0010, 1'b0, 1'b0); // 2 % 5 = 2
  run_test(4'b1000, 4'b0011, 6'b001101, 4'b0010, 1'b0, 1'b0); // 8 % 3 = 2

  // when Sel is 6'b010100 which indicates Parity_Checker( A ) 
  run_test(4'b0000, 4'b1000, 6'b010100, 4'b0000, 1'b0, 1'b0); // A = 0000 → 0 ones → even
  run_test(4'b0001, 4'b1000, 6'b010100, 4'b0001, 1'b0, 1'b0); // A = 0001 → 1 one  → odd
  run_test(4'b0011, 4'b1000, 6'b010100, 4'b0000, 1'b0, 1'b0); // A = 0011 → 2 ones → even
  run_test(4'b0101, 4'b1000, 6'b010100, 4'b0000, 1'b0, 1'b0); // A = 0101 → 2 ones → even
  run_test(4'b0110, 4'b1000, 6'b010100, 4'b0000, 1'b0, 1'b0); // A = 0110 → 2 ones → even
  run_test(4'b0111, 4'b1000, 6'b010100, 4'b0001, 1'b0, 1'b0); // A = 0111 → 3 ones → odd
  run_test(4'b1000, 4'b1000, 6'b010100, 4'b0001, 1'b0, 1'b0); // A = 1000 → 1 one  → odd
  run_test(4'b1111, 4'b1000, 6'b010100, 4'b0000, 1'b0, 1'b0); // A = 1111 → 4 ones → even
  run_test(4'b1010, 4'b1000, 6'b010100, 4'b0000, 1'b0, 1'b0); // A = 1010 → 2 ones → even

  // when Sel is 6'b010101 which indicates Parity_Checker( B ) 
  run_test(4'b0101, 4'b0000, 6'b010101, 4'b0000, 1'b0, 1'b0); // B = 0000 → 0 ones → even
  run_test(4'b1100, 4'b0001, 6'b010101, 4'b0001, 1'b0, 1'b0); // B = 0001 → 1 one  → odd
  run_test(4'b0001, 4'b0011, 6'b010101, 4'b0000, 1'b0, 1'b0); // B = 0011 → 2 ones → even
  run_test(4'b0011, 4'b0101, 6'b010101, 4'b0000, 1'b0, 1'b0); // B = 0101 → 2 ones → even
  run_test(4'b1010, 4'b0110, 6'b010101, 4'b0000, 1'b0, 1'b0); // B = 0110 → 2 ones → even
  run_test(4'b1101, 4'b0111, 6'b010101, 4'b0001, 1'b0, 1'b0); // B = 0111 → 3 ones → odd
  run_test(4'b0001, 4'b1000, 6'b010101, 4'b0001, 1'b0, 1'b0); // B = 1000 → 1 one  → odd
  run_test(4'b0010, 4'b1111, 6'b010101, 4'b0000, 1'b0, 1'b0); // B = 1111 → 4 ones → even
  run_test(4'b1000, 4'b1010, 6'b010101, 4'b0000, 1'b0, 1'b0); // B = 1010 → 2 ones → even

  // when Sel is 6'b001010 which indicates Arithmetic Shift Right ( A ) 
  run_test(4'b0101, 4'b1000, 6'b001010, 4'b0010, 1'b0, 1'b0); // 0101 >> 1 = 0010
  run_test(4'b1100, 4'b1000, 6'b001010, 4'b1110, 1'b0, 1'b0); // 1100 >> 1 = 1110
  run_test(4'b0001, 4'b1000, 6'b001010, 4'b0000, 1'b0, 1'b0); // 0001 >> 1 = 0000
  run_test(4'b0011, 4'b1000, 6'b001010, 4'b0001, 1'b0, 1'b0); // 0011 >> 1 = 0001
  run_test(4'b1010, 4'b1000, 6'b001010, 4'b1101, 1'b0, 1'b0); // 1010 >> 1 = 1101
  run_test(4'b1101, 4'b1000, 6'b001010, 4'b1110, 1'b0, 1'b0); // 1101 >> 1 = 1110
  run_test(4'b0001, 4'b1000, 6'b001010, 4'b0000, 1'b0, 1'b0); // 0001 >> 1 = 0000
  run_test(4'b0010, 4'b1000, 6'b001010, 4'b0001, 1'b0, 1'b0); // 0010 >> 1 = 0001
  run_test(4'b1000, 4'b1000, 6'b001010, 4'b1100, 1'b0, 1'b0); // 1000 >> 1 = 1100

  // when Sel is 6'b001111 which indicates Arithmetic Shift Left ( A ) 
  run_test(4'b0101, 4'b1000, 6'b001111, 4'b1010, 1'b0, 1'b0); // 0101 << 1 = 1010
  run_test(4'b1100, 4'b1000, 6'b001111, 4'b1000, 1'b0, 1'b0); // 1100 << 1 = 1000
  run_test(4'b0001, 4'b1000, 6'b001111, 4'b0010, 1'b0, 1'b0); // 0001 << 1 = 0010
  run_test(4'b0011, 4'b1000, 6'b001111, 4'b0110, 1'b0, 1'b0); // 0011 << 1 = 0110
  run_test(4'b1010, 4'b1000, 6'b001111, 4'b0100, 1'b0, 1'b0); // 1010 << 1 = 0100
  run_test(4'b1101, 4'b1000, 6'b001111, 4'b1010, 1'b0, 1'b0); // 1101 << 1 = 1010
  run_test(4'b0001, 4'b1000, 6'b001111, 4'b0010, 1'b0, 1'b0); // 0001 << 1 = 0010
  run_test(4'b0010, 4'b1000, 6'b001111, 4'b0100, 1'b0, 1'b0); // 0010 << 1 = 0100
  run_test(4'b1000, 4'b1000, 6'b001111, 4'b0000, 1'b0, 1'b0); // 1000 << 1 = 0000 

  // when Sel is 6'b011011 which indicates Arithmetic Shift Right ( B ) 
  run_test(4'b0101, 4'b0001, 6'b011011, 4'b0000, 1'b0, 1'b0); // 0001 >>> 1 = 0000
  run_test(4'b1100, 4'b0010, 6'b011011, 4'b0001, 1'b0, 1'b0); // 0010 >>> 1 = 0001
  run_test(4'b0001, 4'b0100, 6'b011011, 4'b0010, 1'b0, 1'b0); // 0100 >>> 1 = 0010
  run_test(4'b0011, 4'b0110, 6'b011011, 4'b0011, 1'b0, 1'b0); // 0110 >>> 1 = 0011
  run_test(4'b1010, 4'b1000, 6'b011011, 4'b1100, 1'b0, 1'b0); // 1000 >>> 1 = 1100 
  run_test(4'b1101, 4'b1010, 6'b011011, 4'b1101, 1'b0, 1'b0); // 1010 >>> 1 = 1101
  run_test(4'b0001, 4'b1100, 6'b011011, 4'b1110, 1'b0, 1'b0); // 1100 >>> 1 = 1110
  run_test(4'b0010, 4'b1110, 6'b011011, 4'b1111, 1'b0, 1'b0); // 1110 >>> 1 = 1111
  run_test(4'b1000, 4'b1111, 6'b011011, 4'b1111, 1'b0, 1'b0); // 1111 >>> 1 = 1111


  // when Sel is 6'b011111 which indicates Arithmetic Shift Left ( B )
  run_test(4'b0101, 4'b0001, 6'b011111, 4'b0010, 1'b0, 1'b0); // 0001 << 1 = 0010
  run_test(4'b1100, 4'b0010, 6'b011111, 4'b0100, 1'b0, 1'b0); // 0010 << 1 = 0100
  run_test(4'b0001, 4'b0011, 6'b011111, 4'b0110, 1'b0, 1'b0); // 0011 << 1 = 0110
  run_test(4'b0011, 4'b0100, 6'b011111, 4'b1000, 1'b0, 1'b0); // 0100 << 1 = 1000
  run_test(4'b1010, 4'b0101, 6'b011111, 4'b1010, 1'b0, 1'b0); // 0101 << 1 = 1010
  run_test(4'b1101, 4'b0110, 6'b011111, 4'b1100, 1'b0, 1'b0); // 0110 << 1 = 1100
  run_test(4'b0001, 4'b0111, 6'b011111, 4'b1110, 1'b0, 1'b0); // 0111 << 1 = 1110
  run_test(4'b0010, 4'b1000, 6'b011111, 4'b0000, 1'b0, 1'b0); // 1000 << 1 = 0000 
  run_test(4'b1000, 4'b1111, 6'b011111, 4'b1110, 1'b0, 1'b0); // 1111 << 1 = 1110 

  // when Sel is 6'b010000 which indicates Reverse ( A )
  run_test(4'b0101, 4'b1000, 6'b010000, 4'b1010, 1'b0, 1'b0); // A = 0101 -> 1010
  run_test(4'b1100, 4'b1000, 6'b010000, 4'b0011, 1'b0, 1'b0); // A = 1100 -> 0011
  run_test(4'b0001, 4'b1000, 6'b010000, 4'b1000, 1'b0, 1'b0); // A = 0001 -> 1000
  run_test(4'b0011, 4'b1000, 6'b010000, 4'b1100, 1'b0, 1'b0); // A = 0011 -> 1100
  run_test(4'b1010, 4'b1000, 6'b010000, 4'b0101, 1'b0, 1'b0); // A = 1010 -> 0101
  run_test(4'b1101, 4'b1000, 6'b010000, 4'b1011, 1'b0, 1'b0); // A = 1101 -> 1011
  run_test(4'b0110, 4'b1000, 6'b010000, 4'b0110, 1'b0, 1'b0); // A = 0110 -> 0110
  run_test(4'b1111, 4'b1000, 6'b010000, 4'b1111, 1'b0, 1'b0); // A = 1111 -> 1111
  run_test(4'b1000, 4'b1000, 6'b010000, 4'b0001, 1'b0, 1'b0); // A = 1000 -> 0001

  // when Sel is 6'b010001 which indicates Reverse ( B )
  run_test(4'b0101, 4'b1000, 6'b010001, 4'b0001, 1'b0, 1'b0); // B = 1000 -> 0001
  run_test(4'b1100, 4'b0001, 6'b010001, 4'b1000, 1'b0, 1'b0); // B = 0001 -> 1000
  run_test(4'b0001, 4'b0011, 6'b010001, 4'b1100, 1'b0, 1'b0); // B = 0011 -> 1100
  run_test(4'b0011, 4'b0101, 6'b010001, 4'b1010, 1'b0, 1'b0); // B = 0101 -> 1010
  run_test(4'b1010, 4'b1110, 6'b010001, 4'b0111, 1'b0, 1'b0); // B = 1110 -> 0111
  run_test(4'b1101, 4'b1010, 6'b010001, 4'b0101, 1'b0, 1'b0); // B = 1010 -> 0101
  run_test(4'b0001, 4'b1001, 6'b010001, 4'b1001, 1'b0, 1'b0); // B = 1001 -> 1001
  run_test(4'b0010, 4'b1111, 6'b010001, 4'b1111, 1'b0, 1'b0); // B = 1111 -> 1111
  run_test(4'b1000, 4'b0110, 6'b010001, 4'b0110, 1'b0, 1'b0); // B = 0110 -> 0110

  // when Sel is 6'b011100 which indicates Increment ( A )
  run_test(4'b0101, 4'b1000, 6'b011100, 4'b0110, 1'b0, 1'b0); // 0101 + 1 = 0110
  run_test(4'b1100, 4'b1000, 6'b011100, 4'b1101, 1'b0, 1'b0); // 1100 + 1 = 1101
  run_test(4'b0001, 4'b1000, 6'b011100, 4'b0010, 1'b0, 1'b0); // 0001 + 1 = 0010
  run_test(4'b0011, 4'b1000, 6'b011100, 4'b0100, 1'b0, 1'b0); // 0011 + 1 = 0100
  run_test(4'b1010, 4'b1000, 6'b011100, 4'b1011, 1'b0, 1'b0); // 1010 + 1 = 1011
  run_test(4'b1101, 4'b1000, 6'b011100, 4'b1110, 1'b0, 1'b0); // 1101 + 1 = 1110
  run_test(4'b1111, 4'b1000, 6'b011100, 4'b0000, 1'b1, 1'b0); // 1111 + 1 = 0000, Carry_Out = 1
  run_test(4'b0000, 4'b1000, 6'b011100, 4'b0001, 1'b0, 1'b0); // 0000 + 1 = 0001
  run_test(4'b0111, 4'b1000, 6'b011100, 4'b1000, 1'b0, 1'b0); // 0111 + 1 = 1000

  // when Sel is 6'b011101 which indicates Increment ( B )
  run_test(4'b0101, 4'b1000, 6'b011101, 4'b1001, 1'b0, 1'b0); // 1000 + 1 = 1001
  run_test(4'b1100, 4'b0111, 6'b011101, 4'b1000, 1'b0, 1'b0); // 0111 + 1 = 1000
  run_test(4'b0001, 4'b0000, 6'b011101, 4'b0001, 1'b0, 1'b0); // 0000 + 1 = 0001
  run_test(4'b0011, 4'b0001, 6'b011101, 4'b0010, 1'b0, 1'b0); // 0001 + 1 = 0010
  run_test(4'b1010, 4'b0010, 6'b011101, 4'b0011, 1'b0, 1'b0); // 0010 + 1 = 0011
  run_test(4'b1101, 4'b1110, 6'b011101, 4'b1111, 1'b0, 1'b0); // 1110 + 1 = 1111
  run_test(4'b0001, 4'b1001, 6'b011101, 4'b1010, 1'b0, 1'b0); // 1001 + 1 = 1010
  run_test(4'b0010, 4'b1111, 6'b011101, 4'b0000, 1'b1, 1'b0); // 1111 + 1 = 0000, Carry_Out = 1
  run_test(4'b1000, 4'b0111, 6'b011101, 4'b1000, 1'b0, 1'b0); // 0111 + 1 = 1000

  // when Sel is 6'b011000 which indicates Decrement(A)
  run_test(4'b0101, 4'b1000, 6'b011000, 4'b0100, 1'b0, 1'b0); // 0101 - 1 = 0100
  run_test(4'b1100, 4'b1000, 6'b011000, 4'b1011, 1'b0, 1'b0); // 1100 - 1 = 1011
  run_test(4'b0001, 4'b1000, 6'b011000, 4'b0000, 1'b0, 1'b0); // 0001 - 1 = 0000
  run_test(4'b0011, 4'b1000, 6'b011000, 4'b0010, 1'b0, 1'b0); // 0011 - 1 = 0010
  run_test(4'b1010, 4'b1000, 6'b011000, 4'b1001, 1'b0, 1'b0); // 1010 - 1 = 1001
  run_test(4'b1101, 4'b1000, 6'b011000, 4'b1100, 1'b0, 1'b0); // 1101 - 1 = 1100
  run_test(4'b0111, 4'b1000, 6'b011000, 4'b0110, 1'b0, 1'b0); // 0111 - 1 = 0110
  run_test(4'b0010, 4'b1000, 6'b011000, 4'b0001, 1'b0, 1'b0); // 0010 - 1 = 0001
  run_test(4'b1000, 4'b1000, 6'b011000, 4'b0111, 1'b0, 1'b0); // 1000 - 1 = 0111
  run_test(4'b0000, 4'b1000, 6'b011000, 4'b0001, 1'b0, 1'b1); // 0000 - 1 = 0001 (but Negative) 

  // when Sel is 6'b011001 which indicates Decrement ( B ) 
  run_test(4'b0000, 4'b0101, 6'b011001, 4'b0100, 1'b0, 1'b0); // 0101 - 1 = 0100
  run_test(4'b0000, 4'b1100, 6'b011001, 4'b1011, 1'b0, 1'b0); // 1100 - 1 = 1011
  run_test(4'b0000, 4'b0001, 6'b011001, 4'b0000, 1'b0, 1'b0); // 0001 - 1 = 0000
  run_test(4'b0000, 4'b0011, 6'b011001, 4'b0010, 1'b0, 1'b0); // 0011 - 1 = 0010
  run_test(4'b0000, 4'b1010, 6'b011001, 4'b1001, 1'b0, 1'b0); // 1010 - 1 = 1001
  run_test(4'b0000, 4'b1101, 6'b011001, 4'b1100, 1'b0, 1'b0); // 1101 - 1 = 1100
  run_test(4'b0000, 4'b0111, 6'b011001, 4'b0110, 1'b0, 1'b0); // 0111 - 1 = 0110
  run_test(4'b0000, 4'b0010, 6'b011001, 4'b0001, 1'b0, 1'b0); // 0010 - 1 = 0001
  run_test(4'b0000, 4'b1000, 6'b011001, 4'b0111, 1'b0, 1'b0); // 1000 - 1 = 0111
  run_test(4'b0000, 4'b0000, 6'b011001, 4'b0001, 1'b0, 1'b1); // 0000 - 1 = 0001 (but Negative)


// --------------------------------------------------------------------------------------------------------------------------------------------

// Logic & Logical Shift Operations

  // when Sel is 6'b100000 which indicates A & B
  run_test(4'b0101, 4'b1000, 6'b100000, 4'b0000, 1'b0, 1'b0); // 0101 & 1000 = 0000
  run_test(4'b1100, 4'b1000, 6'b100000, 4'b1000, 1'b0, 1'b0); // 1100 & 1000 = 1000
  run_test(4'b0001, 4'b1000, 6'b100000, 4'b0000, 1'b0, 1'b0); // 0001 & 1000 = 0000
  run_test(4'b0011, 4'b1000, 6'b100000, 4'b0000, 1'b0, 1'b0); // 0011 & 1000 = 0000
  run_test(4'b1010, 4'b1000, 6'b100000, 4'b1000, 1'b0, 1'b0); // 1010 & 1000 = 1000
  run_test(4'b1101, 4'b1000, 6'b100000, 4'b1000, 1'b0, 1'b0); // 1101 & 1000 = 1000
  run_test(4'b0001, 4'b1000, 6'b100000, 4'b0000, 1'b0, 1'b0); // 0001 & 1000 = 0000
  run_test(4'b0010, 4'b1000, 6'b100000, 4'b0000, 1'b0, 1'b0); // 0010 & 1000 = 0000
  run_test(4'b1000, 4'b1000, 6'b100000, 4'b1000, 1'b0, 1'b0); // 1000 & 1000 = 1000

  // when Sel is 6'b100001 which indicates A | B 
  run_test(4'b0101, 4'b1000, 6'b100001, 4'b1101, 1'b0, 1'b0); // 0101 | 1000 = 1101
  run_test(4'b1100, 4'b1000, 6'b100001, 4'b1100, 1'b0, 1'b0); // 1100 | 1000 = 1100
  run_test(4'b0001, 4'b1000, 6'b100001, 4'b1001, 1'b0, 1'b0); // 0001 | 1000 = 1001
  run_test(4'b0011, 4'b1000, 6'b100001, 4'b1011, 1'b0, 1'b0); // 0011 | 1000 = 1011
  run_test(4'b1010, 4'b1000, 6'b100001, 4'b1010, 1'b0, 1'b0); // 1010 | 1000 = 1010
  run_test(4'b1101, 4'b1000, 6'b100001, 4'b1101, 1'b0, 1'b0); // 1101 | 1000 = 1101
  run_test(4'b0001, 4'b1000, 6'b100001, 4'b1001, 1'b0, 1'b0); // 0001 | 1000 = 1001
  run_test(4'b0010, 4'b1000, 6'b100001, 4'b1010, 1'b0, 1'b0); // 0010 | 1000 = 1010
  run_test(4'b1000, 4'b1000, 6'b100001, 4'b1000, 1'b0, 1'b0); // 1000 | 1000 = 1000

  // when Sel is 6'b100010 which indicates A ^ B 
  run_test(4'b0101, 4'b1000, 6'b100010, 4'b1101, 1'b0, 1'b0); // 0101 ^ 1000 = 1101
  run_test(4'b1100, 4'b1000, 6'b100010, 4'b0100, 1'b0, 1'b0); // 1100 ^ 1000 = 0100
  run_test(4'b0001, 4'b1000, 6'b100010, 4'b1001, 1'b0, 1'b0); // 0001 ^ 1000 = 1001
  run_test(4'b0011, 4'b1000, 6'b100010, 4'b1011, 1'b0, 1'b0); // 0011 ^ 1000 = 1011
  run_test(4'b1010, 4'b1000, 6'b100010, 4'b0010, 1'b0, 1'b0); // 1010 ^ 1000 = 0010
  run_test(4'b1101, 4'b1000, 6'b100010, 4'b0101, 1'b0, 1'b0); // 1101 ^ 1000 = 0101
  run_test(4'b0001, 4'b1000, 6'b100010, 4'b1001, 1'b0, 1'b0); // 0001 ^ 1000 = 1001
  run_test(4'b0010, 4'b1000, 6'b100010, 4'b1010, 1'b0, 1'b0); // 0010 ^ 1000 = 1010
  run_test(4'b1000, 4'b1000, 6'b100010, 4'b0000, 1'b0, 1'b0); // 1000 ^ 1000 = 0000

  // when Sel is 6'b100011 which indicates ~(A ^ B)
  run_test(4'b0101, 4'b1000, 6'b100011, 4'b0010, 1'b0, 1'b0); // ~(0101 ^ 1000) = ~(1101) = 0010
  run_test(4'b1100, 4'b1000, 6'b100011, 4'b1011, 1'b0, 1'b0); // ~(1100 ^ 1000) = ~(0100) = 1011
  run_test(4'b0001, 4'b1000, 6'b100011, 4'b0110, 1'b0, 1'b0); // ~(0001 ^ 1000) = ~(1001) = 0110
  run_test(4'b0011, 4'b1000, 6'b100011, 4'b0100, 1'b0, 1'b0); // ~(0011 ^ 1000) = ~(1011) = 0100
  run_test(4'b1010, 4'b1000, 6'b100011, 4'b1101, 1'b0, 1'b0); // ~(1010 ^ 1000) = ~(0010) = 1101
  run_test(4'b1101, 4'b1000, 6'b100011, 4'b1100, 1'b0, 1'b0); // ~(1101 ^ 1000) = ~(0101) = 1010
  run_test(4'b0001, 4'b1000, 6'b100011, 4'b0110, 1'b0, 1'b0); // ~(0001 ^ 1000) = ~(1001) = 0110
  run_test(4'b0010, 4'b1000, 6'b100011, 4'b0101, 1'b0, 1'b0); // ~(0010 ^ 1000) = ~(1010) = 0101
  run_test(4'b1000, 4'b1000, 6'b100011, 4'b1111, 1'b0, 1'b0); // ~(1000 ^ 1000) = ~(0000) = 1111

  // when Sel is 6'b101100 which indicates ~(A & B)
  run_test(4'b0101, 4'b1000, 6'b101100, 4'b1111, 1'b0, 1'b0); // ~(0101 & 1000) = ~(0000) = 1111
  run_test(4'b1100, 4'b1000, 6'b101100, 4'b1011, 1'b0, 1'b0); // ~(1100 & 1000) = ~(1000) = 0111
  run_test(4'b0001, 4'b1000, 6'b101100, 4'b1111, 1'b0, 1'b0); // ~(0001 & 1000) = ~(0000) = 1111
  run_test(4'b0011, 4'b1000, 6'b101100, 4'b1111, 1'b0, 1'b0); // ~(0011 & 1000) = ~(0000) = 1111
  run_test(4'b1010, 4'b1000, 6'b101100, 4'b1111, 1'b0, 1'b0); // ~(1010 & 1000) = ~(1000) = 0111
  run_test(4'b1101, 4'b1000, 6'b101100, 4'b0111, 1'b0, 1'b0); // ~(1101 & 1000) = ~(1000) = 0111
  run_test(4'b0001, 4'b1000, 6'b101100, 4'b1111, 1'b0, 1'b0); // ~(0001 & 1000) = ~(0000) = 1111
  run_test(4'b0010, 4'b1000, 6'b101100, 4'b1111, 1'b0, 1'b0); // ~(0010 & 1000) = ~(0000) = 1111
  run_test(4'b1000, 4'b1000, 6'b101100, 4'b0111, 1'b0, 1'b0); // ~(1000 & 1000) = ~(1000) = 0111

  // when Sel is 6'b101101 which indicates ~(A | B)
  run_test(4'b0101, 4'b1000, 6'b101101, 4'b0010, 1'b0, 1'b0); // ~(0101 | 1000) = ~(1101) = 0010
  run_test(4'b1100, 4'b1000, 6'b101101, 4'b0011, 1'b0, 1'b0); // ~(1100 | 1000) = ~(1100) = 0011
  run_test(4'b0001, 4'b1000, 6'b101101, 4'b0110, 1'b0, 1'b0); // ~(0001 | 1000) = ~(1001) = 0110
  run_test(4'b0011, 4'b1000, 6'b101101, 4'b0100, 1'b0, 1'b0); // ~(0011 | 1000) = ~(1011) = 0100
  run_test(4'b1010, 4'b1000, 6'b101101, 4'b0101, 1'b0, 1'b0); // ~(1010 | 1000) = ~(1010) = 0101
  run_test(4'b1101, 4'b1000, 6'b101101, 4'b0000, 1'b0, 1'b0); // ~(1101 | 1000) = ~(1101) = 0010
  run_test(4'b0001, 4'b1000, 6'b101101, 4'b0110, 1'b0, 1'b0); // ~(0001 | 1000) = ~(1001) = 0110
  run_test(4'b0010, 4'b1000, 6'b101101, 4'b0101, 1'b0, 1'b0); // ~(0010 | 1000) = ~(1010) = 0101
  run_test(4'b1000, 4'b1000, 6'b101101, 4'b0111, 1'b0, 1'b0); // ~(1000 | 1000) = ~(1000) = 0111

  // when Sel is 6'b101110 which indicates ~( A )
  run_test(4'b0101, 4'b1000, 6'b101110, 4'b1010, 1'b0, 1'b0); // ~0101 = 1010
  run_test(4'b1100, 4'b1000, 6'b101110, 4'b0011, 1'b0, 1'b0); // ~1100 = 0011
  run_test(4'b0001, 4'b1000, 6'b101110, 4'b1110, 1'b0, 1'b0); // ~0001 = 1110
  run_test(4'b0011, 4'b1000, 6'b101110, 4'b1100, 1'b0, 1'b0); // ~0011 = 1100
  run_test(4'b1010, 4'b1000, 6'b101110, 4'b0101, 1'b0, 1'b0); // ~1010 = 0101
  run_test(4'b1101, 4'b1000, 6'b101110, 4'b0010, 1'b0, 1'b0); // ~1101 = 0010
  run_test(4'b0001, 4'b1000, 6'b101110, 4'b1110, 1'b0, 1'b0); // ~0001 = 1110
  run_test(4'b0010, 4'b1000, 6'b101110, 4'b1101, 1'b0, 1'b0); // ~0010 = 1101
  run_test(4'b1000, 4'b1000, 6'b101110, 4'b0111, 1'b0, 1'b0); // ~1000 = 0111

  // when Sel is 6'b101111 which indicates ~( B )
  run_test(4'b0101, 4'b1000, 6'b101111, 4'b0111, 1'b0, 1'b0); // ~1000 = 0111
  run_test(4'b1100, 4'b1000, 6'b101111, 4'b0111, 1'b0, 1'b0); // ~1000 = 0111
  run_test(4'b0001, 4'b1000, 6'b101111, 4'b0111, 1'b0, 1'b0); // ~1000 = 0111
  run_test(4'b0011, 4'b1000, 6'b101111, 4'b0111, 1'b0, 1'b0); // ~1000 = 0111
  run_test(4'b1010, 4'b1000, 6'b101111, 4'b0111, 1'b0, 1'b0); // ~1000 = 0111
  run_test(4'b1101, 4'b1000, 6'b101111, 4'b0111, 1'b0, 1'b0); // ~1000 = 0111
  run_test(4'b0001, 4'b1000, 6'b101111, 4'b0111, 1'b0, 1'b0); // ~1000 = 0111
  run_test(4'b0010, 4'b1000, 6'b101111, 4'b0111, 1'b0, 1'b0); // ~1000 = 0111
  run_test(4'b1000, 4'b1000, 6'b101111, 4'b0111, 1'b0, 1'b0); // ~1000 = 0111

  // when Sel is 6'b110000 which indicates ( A )
  run_test(4'b0101, 4'b1000, 6'b110000, 4'b0101, 1'b0, 1'b0); // A = 0101
  run_test(4'b1100, 4'b1000, 6'b110000, 4'b1100, 1'b0, 1'b0); // A = 1100
  run_test(4'b0001, 4'b1000, 6'b110000, 4'b0001, 1'b0, 1'b0); // A = 0001
  run_test(4'b0011, 4'b1000, 6'b110000, 4'b0011, 1'b0, 1'b0); // A = 0011
  run_test(4'b1010, 4'b1000, 6'b110000, 4'b1010, 1'b0, 1'b0); // A = 1010
  run_test(4'b1101, 4'b1000, 6'b110000, 4'b1101, 1'b0, 1'b0); // A = 1101
  run_test(4'b0001, 4'b1000, 6'b110000, 4'b0001, 1'b0, 1'b0); // A = 0001
  run_test(4'b0010, 4'b1000, 6'b110000, 4'b0010, 1'b0, 1'b0); // A = 0010
  run_test(4'b1000, 4'b1000, 6'b110000, 4'b1000, 1'b0, 1'b0); // A = 1000

  // when Sel is 6'b110001 which indicates ( B ) 
  run_test(4'b0000, 4'b0001, 6'b110001, 4'b0001, 1'b0, 1'b0); // B = 0001
  run_test(4'b0000, 4'b0010, 6'b110001, 4'b0010, 1'b0, 1'b0); // B = 0010
  run_test(4'b0000, 4'b0011, 6'b110001, 4'b0011, 1'b0, 1'b0); // B = 0011
  run_test(4'b0000, 4'b0100, 6'b110001, 4'b0100, 1'b0, 1'b0); // B = 0100
  run_test(4'b0000, 4'b0101, 6'b110001, 4'b0101, 1'b0, 1'b0); // B = 0101
  run_test(4'b0000, 4'b0110, 6'b110001, 4'b0110, 1'b0, 1'b0); // B = 0110
  run_test(4'b0000, 4'b0111, 6'b110001, 4'b0111, 1'b0, 1'b0); // B = 0111
  run_test(4'b0000, 4'b1000, 6'b110001, 4'b1000, 1'b0, 1'b0); // B = 1000
  run_test(4'b0000, 4'b1111, 6'b110001, 4'b1111, 1'b0, 1'b0); // B = 1111

  // when Sel is 6'b110010 which indicates if ( A == B ) → 0001 else → 0000 
  run_test(4'b0101, 4'b1000, 6'b110010, 4'b0000, 1'b0, 1'b0); // A ≠ B → 0000
  run_test(4'b1100, 4'b1000, 6'b110010, 4'b0000, 1'b0, 1'b0); // A ≠ B → 0000
  run_test(4'b0001, 4'b1000, 6'b110010, 4'b0000, 1'b0, 1'b0); // A ≠ B → 0000
  run_test(4'b0011, 4'b1000, 6'b110010, 4'b0000, 1'b0, 1'b0); // A ≠ B → 0000
  run_test(4'b1010, 4'b1000, 6'b110010, 4'b0000, 1'b0, 1'b0); // A ≠ B → 0000
  run_test(4'b1101, 4'b1000, 6'b110010, 4'b0000, 1'b0, 1'b0); // A ≠ B → 0000
  run_test(4'b0001, 4'b1000, 6'b110010, 4'b0000, 1'b0, 1'b0); // A ≠ B → 0000
  run_test(4'b0010, 4'b1000, 6'b110010, 4'b0000, 1'b0, 1'b0); // A ≠ B → 0000
  run_test(4'b1000, 4'b1000, 6'b110010, 4'b0001, 1'b0, 1'b0); // A == B → 0001
  run_test(4'b0000, 4'b0000, 6'b110010, 4'b0001, 1'b0, 1'b0); // A == B → 0001
  run_test(4'b1111, 4'b1111, 6'b110010, 4'b0001, 1'b0, 1'b0); // A == B → 0001
  run_test(4'b1010, 4'b1010, 6'b110010, 4'b0001, 1'b0, 1'b0); // A == B → 0001
  run_test(4'b0101, 4'b0101, 6'b110010, 4'b0001, 1'b0, 1'b0); // A == B → 0001

  // when Sel is 6'b110011 which indicates if ( A < B ) output ==> 4'b0001 and otherwise 4'b0000 
  run_test(4'b0101, 4'b1000, 6'b110011, 4'b0001, 1'b0, 1'b0); // 5 < 8 → 0001
  run_test(4'b1100, 4'b1000, 6'b110011, 4'b0000, 1'b0, 1'b0); // 12 > 8 → 0000
  run_test(4'b0001, 4'b1000, 6'b110011, 4'b0001, 1'b0, 1'b0); // 1 < 8 → 0001
  run_test(4'b0011, 4'b1000, 6'b110011, 4'b0001, 1'b0, 1'b0); // 3 < 8 → 0001
  run_test(4'b1010, 4'b1000, 6'b110011, 4'b0000, 1'b0, 1'b0); // 10 > 8 → 0000
  run_test(4'b1101, 4'b1000, 6'b110011, 4'b0000, 1'b0, 1'b0); // 13 > 8 → 0000
  run_test(4'b0001, 4'b1000, 6'b110011, 4'b0001, 1'b0, 1'b0); // 1 < 8 → 0001
  run_test(4'b0010, 4'b1000, 6'b110011, 4'b0001, 1'b0, 1'b0); // 2 < 8 → 0001
  run_test(4'b1000, 4'b1000, 6'b110011, 4'b0000, 1'b0, 1'b0); // 8 == 8 → 0000

  // when Sel is 6'b111000 which indicates Logic Shift Right ( A )
  run_test(4'b0101, 4'b1000, 6'b111000, 4'b0010, 1'b0, 1'b0); // 0101 >> 1 = 0010
  run_test(4'b1100, 4'b1000, 6'b111000, 4'b0110, 1'b0, 1'b0); // 1100 >> 1 = 0110
  run_test(4'b0001, 4'b1000, 6'b111000, 4'b0000, 1'b0, 1'b0); // 0001 >> 1 = 0000
  run_test(4'b0011, 4'b1000, 6'b111000, 4'b0001, 1'b0, 1'b0); // 0011 >> 1 = 0001
  run_test(4'b1010, 4'b1000, 6'b111000, 4'b0101, 1'b0, 1'b0); // 1010 >> 1 = 0101
  run_test(4'b1101, 4'b1000, 6'b111000, 4'b0110, 1'b0, 1'b0); // 1101 >> 1 = 0110
  run_test(4'b0001, 4'b1000, 6'b111000, 4'b0000, 1'b0, 1'b0); // 0001 >> 1 = 0000
  run_test(4'b0010, 4'b1000, 6'b111000, 4'b0001, 1'b0, 1'b0); // 0010 >> 1 = 0001
  run_test(4'b1000, 4'b1000, 6'b111000, 4'b0100, 1'b0, 1'b0); // 1000 >> 1 = 0100

  // when Sel is 6'b111001 which indicates Logic Shift Left ( A )
  run_test(4'b0101, 4'b1000, 6'b111001, 4'b1010, 1'b0, 1'b0); // 0101 << 1 = 1010
  run_test(4'b1100, 4'b1000, 6'b111001, 4'b1000, 1'b0, 1'b0); // 1100 << 1 = 1000
  run_test(4'b0001, 4'b1000, 6'b111001, 4'b0010, 1'b0, 1'b0); // 0001 << 1 = 0010
  run_test(4'b0011, 4'b1000, 6'b111001, 4'b0110, 1'b0, 1'b0); // 0011 << 1 = 0110
  run_test(4'b1010, 4'b1000, 6'b111001, 4'b0100, 1'b0, 1'b0); // 1010 << 1 = 0100
  run_test(4'b1101, 4'b1000, 6'b111001, 4'b1010, 1'b0, 1'b0); // 1101 << 1 = 1010
  run_test(4'b0001, 4'b1000, 6'b111001, 4'b0010, 1'b0, 1'b0); // 0001 << 1 = 0010
  run_test(4'b0010, 4'b1000, 6'b111001, 4'b0100, 1'b0, 1'b0); // 0010 << 1 = 0100
  run_test(4'b1000, 4'b1000, 6'b111001, 4'b0000, 1'b0, 1'b0); // 1000 << 1 = 0000 (MSB dropped)

  // when Sel is 6'b111010 which indicates Logic Shift Right ( B )
  run_test(4'b0101, 4'b1000, 6'b111010, 4'b0100, 1'b0, 1'b0); // 1000 >> 1 = 0100
  run_test(4'b1100, 4'b0100, 6'b111010, 4'b0010, 1'b0, 1'b0); // 0100 >> 1 = 0010
  run_test(4'b0001, 4'b0001, 6'b111010, 4'b0000, 1'b0, 1'b0); // 0001 >> 1 = 0000
  run_test(4'b0011, 4'b0010, 6'b111010, 4'b0001, 1'b0, 1'b0); // 0010 >> 1 = 0001
  run_test(4'b1010, 4'b1111, 6'b111010, 4'b0111, 1'b0, 1'b0); // 1111 >> 1 = 0111
  run_test(4'b1101, 4'b1010, 6'b111010, 4'b0101, 1'b0, 1'b0); // 1010 >> 1 = 0101
  run_test(4'b0001, 4'b0011, 6'b111010, 4'b0001, 1'b0, 1'b0); // 0011 >> 1 = 0001
  run_test(4'b0010, 4'b0110, 6'b111010, 4'b0011, 1'b0, 1'b0); // 0110 >> 1 = 0011
  run_test(4'b1000, 4'b1001, 6'b111010, 4'b0100, 1'b0, 1'b0); // 1001 >> 1 = 0100

  // when Sel is 6'b111011 which indicates Logic Shift Left ( B )
  run_test(4'b0101, 4'b0001, 6'b111011, 4'b0010, 1'b0, 1'b0); // 0001 << 1 = 0010
  run_test(4'b1100, 4'b0010, 6'b111011, 4'b0100, 1'b0, 1'b0); // 0010 << 1 = 0100
  run_test(4'b0001, 4'b0011, 6'b111011, 4'b0110, 1'b0, 1'b0); // 0011 << 1 = 0110
  run_test(4'b0011, 4'b0100, 6'b111011, 4'b1000, 1'b0, 1'b0); // 0100 << 1 = 1000
  run_test(4'b1010, 4'b1000, 6'b111011, 4'b0000, 1'b0, 1'b0); // 1000 << 1 = 0000 (overflowed bit dropped)
  run_test(4'b1101, 4'b1010, 6'b111011, 4'b0100, 1'b0, 1'b0); // 1010 << 1 = 0100
  run_test(4'b0001, 4'b1100, 6'b111011, 4'b1000, 1'b0, 1'b0); // 1100 << 1 = 1000
  run_test(4'b0010, 4'b1110, 6'b111011, 4'b1100, 1'b0, 1'b0); // 1110 << 1 = 1100
  run_test(4'b1000, 4'b1111, 6'b111011, 4'b1110, 1'b0, 1'b0); // 1111 << 1 = 1110

  // when Sel is 6'b111100 which indicates Rotate Right ( A )
  run_test(4'b0101, 4'b1000, 6'b111100, 4'b1010, 1'b0, 1'b0); // 0101 -> 1010
  run_test(4'b1100, 4'b1000, 6'b111100, 4'b0110, 1'b0, 1'b0); // 1100 -> 0110
  run_test(4'b0001, 4'b1000, 6'b111100, 4'b1000, 1'b0, 1'b0); // 0001 -> 1000
  run_test(4'b0011, 4'b1000, 6'b111100, 4'b1001, 1'b0, 1'b0); // 0011 -> 1001
  run_test(4'b1010, 4'b1000, 6'b111100, 4'b0101, 1'b0, 1'b0); // 1010 -> 0101
  run_test(4'b1101, 4'b1000, 6'b111100, 4'b1110, 1'b0, 1'b0); // 1101 -> 1110
  run_test(4'b0001, 4'b1000, 6'b111100, 4'b1000, 1'b0, 1'b0); // 0001 -> 1000
  run_test(4'b0010, 4'b1000, 6'b111100, 4'b0001, 1'b0, 1'b0); // 0010 -> 0001
  run_test(4'b1000, 4'b1000, 6'b111100, 4'b0100, 1'b0, 1'b0); // 1000 -> 0100

  // when Sel is 6'b111101 which indicates Rotate Left ( A )
  run_test(4'b0101, 4'b1000, 6'b111101, 4'b1010, 1'b0, 1'b0); // 0101 -> 1010
  run_test(4'b1100, 4'b1000, 6'b111101, 4'b1001, 1'b0, 1'b0); // 1100 -> 1001
  run_test(4'b0001, 4'b1000, 6'b111101, 4'b0010, 1'b0, 1'b0); // 0001 -> 0010
  run_test(4'b0011, 4'b1000, 6'b111101, 4'b0110, 1'b0, 1'b0); // 0011 -> 0110
  run_test(4'b1010, 4'b1000, 6'b111101, 4'b0101, 1'b0, 1'b0); // 1010 -> 0101
  run_test(4'b1101, 4'b1000, 6'b111101, 4'b1011, 1'b0, 1'b0); // 1101 -> 1011
  run_test(4'b0001, 4'b1000, 6'b111101, 4'b0010, 1'b0, 1'b0); // 0001 -> 0010
  run_test(4'b0010, 4'b1000, 6'b111101, 4'b0100, 1'b0, 1'b0); // 0010 -> 0100
  run_test(4'b1000, 4'b1000, 6'b111101, 4'b0001, 1'b0, 1'b0); // 1000 -> 0001

  // when Sel is 6'b111110 which indicates Rotate Right ( B )
  run_test(4'b0101, 4'b1000, 6'b111110, 4'b0100, 1'b0, 1'b0); // 1000 -> 0100
  run_test(4'b1100, 4'b0001, 6'b111110, 4'b1000, 1'b0, 1'b0); // 0001 -> 1000
  run_test(4'b0001, 4'b0010, 6'b111110, 4'b0001, 1'b0, 1'b0); // 0010 -> 0001
  run_test(4'b0011, 4'b0011, 6'b111110, 4'b1001, 1'b0, 1'b0); // 0011 -> 1001
  run_test(4'b1010, 4'b0100, 6'b111110, 4'b0010, 1'b0, 1'b0); // 0100 -> 0010
  run_test(4'b1101, 4'b0101, 6'b111110, 4'b1010, 1'b0, 1'b0); // 0101 -> 1010
  run_test(4'b0001, 4'b1111, 6'b111110, 4'b1111, 1'b0, 1'b0); // 1111 -> 1111
  run_test(4'b0010, 4'b1001, 6'b111110, 4'b1100, 1'b0, 1'b0); // 1001 -> 1100
  run_test(4'b1000, 4'b0000, 6'b111110, 4'b0000, 1'b0, 1'b0); // 0000 -> 0000

  // when Sel is 6'b111111 which indicates Rotate Left ( B )
  run_test(4'b0101, 4'b1000, 6'b111111, 4'b0001, 1'b0, 1'b0); // 1000 -> 0001
  run_test(4'b1100, 4'b0001, 6'b111111, 4'b0010, 1'b0, 1'b0); // 0001 -> 0010
  run_test(4'b0001, 4'b0010, 6'b111111, 4'b0100, 1'b0, 1'b0); // 0010 -> 0100
  run_test(4'b0011, 4'b0011, 6'b111111, 4'b0110, 1'b0, 1'b0); // 0011 -> 0110
  run_test(4'b1010, 4'b0100, 6'b111111, 4'b1000, 1'b0, 1'b0); // 0100 -> 1000
  run_test(4'b1101, 4'b0101, 6'b111111, 4'b1010, 1'b0, 1'b0); // 0101 -> 1010
  run_test(4'b0001, 4'b1111, 6'b111111, 4'b1111, 1'b0, 1'b0); // 1111 -> 1111
  run_test(4'b0010, 4'b1001, 6'b111111, 4'b0011, 1'b0, 1'b0); // 1001 -> 0011
  run_test(4'b1000, 4'b0000, 6'b111111, 4'b0000, 1'b0, 1'b0); // 0000 -> 0000

  #Delay;

   if (error_count == 0) begin
      $display("All tests passed successfully!");
    end else begin
      $display("Test completed with %0d errors.", error_count);
    end

    $stop; 
   
  end 

  task run_test(
    input [Width-1:0] a_in,
    input [Width-1:0] b_in,
    input [Width_Sel-1:0] Sel_in,
    input [Output_Width-1:0] expected_out,
    input expected_carry_out,
    input Expected_Sign_Flag
  );
    begin
      A = a_in;
      B = b_in;
      Sel = Sel_in;
      #Delay; 
      if ( (Out !== expected_out) && (carry_out !== expected_carry_out ) && (Expected_Sign_Flag !== Negative_Sign_Flag)) begin
        $display("ERROR at time %0t: A=%b (%0d), B=%b (%0d), Sel=%b (%0d), Expected Out=%b (%0d), Got Out=%b (%0d), Expected Carry=%b (%0d), Got Carry Out=%b (%0d), Expected Sign Flag=%b (%0d)",  
                 $time, A, A, B, B, Sel, Sel, expected_out, expected_out, Out, Out, expected_carry_out, expected_carry_out , carry_out, carry_out , Expected_Sign_Flag , Expected_Sign_Flag , Negative_Sign_Flag , Negative_Sign_Flag);
        error_count = error_count + 1;
      end else begin
        $display("PASS: A=%0d, B=%0d, Sel=%b, Out=%0d", A, B, Sel, Out, carry_out);
      end
    end
  endtask

endmodule 
